module main(
	input sampleInput, 
	output sampleOutput);
	
	assign sampleOutput = sampleInput;

endmodule
